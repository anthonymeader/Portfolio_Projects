-- soc_system_bandpassEQ_ad1939_subsytem.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_bandpassEQ_ad1939_subsytem is
	port (
		ad1939_physical_asdata2     : in  std_logic                     := '0';             --         ad1939_physical.asdata2
		ad1939_physical_dsdata1     : out std_logic;                                        --                        .dsdata1
		ad1939_physical_dbclk       : out std_logic;                                        --                        .dbclk
		ad1939_physical_dlrclk      : out std_logic;                                        --                        .dlrclk
		ad1939_physical_abclk_clk   : in  std_logic                     := '0';             --   ad1939_physical_abclk.clk
		ad1939_physical_alrclk_clk  : in  std_logic                     := '0';             --  ad1939_physical_alrclk.clk
		ad1939_physical_mclk_clk    : in  std_logic                     := '0';             --    ad1939_physical_mclk.clk
		audio_fabric_system_clk_clk : out std_logic;                                        -- audio_fabric_system_clk.clk
		from_line_in_channel        : out std_logic;                                        --            from_line_in.channel
		from_line_in_data           : out std_logic_vector(23 downto 0);                    --                        .data
		from_line_in_valid          : out std_logic;                                        --                        .valid
		subsystem_reset_reset       : in  std_logic                     := '0';             --         subsystem_reset.reset
		to_headphone_out_channel    : in  std_logic                     := '0';             --        to_headphone_out.channel
		to_headphone_out_data       : in  std_logic_vector(23 downto 0) := (others => '0'); --                        .data
		to_headphone_out_valid      : in  std_logic                     := '0'              --                        .valid
	);
end entity soc_system_bandpassEQ_ad1939_subsytem;

architecture rtl of soc_system_bandpassEQ_ad1939_subsytem is
	component ad1939_hps_audio_mini is
		port (
			sys_clk            : in  std_logic                     := 'X';             -- clk
			ad1939_adc_abclk   : in  std_logic                     := 'X';             -- clk
			ad1939_adc_alrclk  : in  std_logic                     := 'X';             -- clk
			sys_reset          : in  std_logic                     := 'X';             -- reset
			ad1939_dac_channel : in  std_logic                     := 'X';             -- channel
			ad1939_dac_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			ad1939_dac_valid   : in  std_logic                     := 'X';             -- valid
			ad1939_adc_channel : out std_logic;                                        -- channel
			ad1939_adc_data    : out std_logic_vector(23 downto 0);                    -- data
			ad1939_adc_valid   : out std_logic;                                        -- valid
			ad1939_adc_asdata2 : in  std_logic                     := 'X';             -- asdata2
			ad1939_dac_dsdata1 : out std_logic;                                        -- dsdata1
			ad1939_dac_dbclk   : out std_logic;                                        -- dbclk
			ad1939_dac_dlrclk  : out std_logic                                         -- dlrclk
		);
	end component ad1939_hps_audio_mini;

	component soc_system_bandpassEQ_ad1939_subsytem_sys_clk_from_ad1939_mclk_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component soc_system_bandpassEQ_ad1939_subsytem_sys_clk_from_ad1939_mclk_pll;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal sys_clk_from_ad1939_mclk_pll_outclk0_clk : std_logic; -- sys_clk_from_ad1939_mclk_pll:outclk_0 -> [audio_fabric_system_clk_clk, AD1939_Audio_Mini:sys_clk, rst_controller:clk]
	signal rst_controller_reset_out_reset           : std_logic; -- rst_controller:reset_out -> AD1939_Audio_Mini:sys_reset

begin

	ad1939_audio_mini : component ad1939_hps_audio_mini
		port map (
			sys_clk            => sys_clk_from_ad1939_mclk_pll_outclk0_clk, --           sys_clk.clk
			ad1939_adc_abclk   => ad1939_physical_abclk_clk,                --         clk_abclk.clk
			ad1939_adc_alrclk  => ad1939_physical_alrclk_clk,               --        clk_alrclk.clk
			sys_reset          => rst_controller_reset_out_reset,           --         sys_reset.reset
			ad1939_dac_channel => to_headphone_out_channel,                 --  to_headphone_out.channel
			ad1939_dac_data    => to_headphone_out_data,                    --                  .data
			ad1939_dac_valid   => to_headphone_out_valid,                   --                  .valid
			ad1939_adc_channel => from_line_in_channel,                     --      from_line_in.channel
			ad1939_adc_data    => from_line_in_data,                        --                  .data
			ad1939_adc_valid   => from_line_in_valid,                       --                  .valid
			ad1939_adc_asdata2 => ad1939_physical_asdata2,                  -- connect_to_AD1939.asdata2
			ad1939_dac_dsdata1 => ad1939_physical_dsdata1,                  --                  .dsdata1
			ad1939_dac_dbclk   => ad1939_physical_dbclk,                    --                  .dbclk
			ad1939_dac_dlrclk  => ad1939_physical_dlrclk                    --                  .dlrclk
		);

	sys_clk_from_ad1939_mclk_pll : component soc_system_bandpassEQ_ad1939_subsytem_sys_clk_from_ad1939_mclk_pll
		port map (
			refclk   => ad1939_physical_mclk_clk,                 --  refclk.clk
			rst      => subsystem_reset_reset,                    --   reset.reset
			outclk_0 => sys_clk_from_ad1939_mclk_pll_outclk0_clk, -- outclk0.clk
			locked   => open                                      -- (terminated)
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => subsystem_reset_reset,                    -- reset_in0.reset
			clk            => sys_clk_from_ad1939_mclk_pll_outclk0_clk, --       clk.clk
			reset_out      => rst_controller_reset_out_reset,           -- reset_out.reset
			reset_req      => open,                                     -- (terminated)
			reset_req_in0  => '0',                                      -- (terminated)
			reset_in1      => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	audio_fabric_system_clk_clk <= sys_clk_from_ad1939_mclk_pll_outclk0_clk;

end architecture rtl; -- of soc_system_bandpassEQ_ad1939_subsytem
